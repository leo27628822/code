
module Comparator( A, B, A_gt_B, A_eq_B, A_lt_B ) ;
// bigger than , equal, less than

input[3:0] A, B;
output A_gt_B, A_eq_B, A_lt_B ;

begin
	
	/* 
	xi = ( A[i] & B[i] ) | ( ~A[i] & ~B[i] ) ;
	assign A_gt_B = ( A[3] & ~B[3] ) | ( x[3] & A[2] & ~B[2] ) | ( x[3] & x[2] & A[1] & ~B[1] ) | ( x[3] & x[2] & x[1] & A[0] & ~B[0] ) ;
	assign A_lt_B = ( ~A[3] & B[3] ) | ( x[3] & ~A[2] & B[2] ) | ( x[3] & x[2] & ~A[1] & B[1] ) | ( x[3] & x[2] & x[1] & ~A[0] & B[0] ) ;
	assign A_eq_B = x[3] & x[2] & x[1] & x[0] ;
	*/
	
	// xi = ( A[] & B[] ) | ( ~A[] & ~B[] ) ;
	assign A_gt_B = ( A[3] & ~B[3] ) | ( ( ( A[3] & B[3] ) | ( ~A[3] & ~B[3] ) ) & A[2] & ~B[2] ) | ( ( ( A[3] & B[3] ) | ( ~A[3] & ~B[3] ) ) & ( ( A[2] & B[2] ) | ( ~A[2] & ~B[2] ) ) & A[1] & ~B[1] ) | ( ( ( A[3] & B[3] ) | ( ~A[3] & ~B[3] ) ) & ( ( A[2] & B[2] ) | ( ~A[2] & ~B[2] ) ) & ( ( A[1] & B[1] ) | ( ~A[1] & ~B[1] ) ) & A[0] & ~B[0] ) ;
	assign A_lt_B = ( ~A[3] & B[3] ) | ( ( ( A[3] & B[3] ) | ( ~A[3] & ~B[3] ) ) & ~A[2] & B[2] ) | ( ( ( A[3] & B[3] ) | ( ~A[3] & ~B[3] ) ) & ( ( A[2] & B[2] ) | ( ~A[2] & ~B[2] ) ) & ~A[1] & B[1] ) | ( ( ( A[3] & B[3] ) | ( ~A[3] & ~B[3] ) ) & ( ( A[2] & B[2] ) | ( ~A[2] & ~B[2] ) ) & ( ( A[1] & B[1] ) | ( ~A[1] & ~B[1] ) ) & ~A[0] & B[0] ) ;
	assign A_eq_B = ( ( A[3] & B[3] ) | ( ~A[3] & ~B[3] ) ) & ( ( A[2] & B[2] ) | ( ~A[2] & ~B[2] ) ) & ( ( A[1] & B[1] ) | ( ~A[1] & ~B[1] ) ) & ( ( A[0] & B[0] ) | ( ~A[0] & ~B[0] ) ) ;

end

endmodule






