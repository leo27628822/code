library verilog;
use verilog.vl_types.all;
entity Counter_10927143 is
    port(
        dout            : out    vl_logic_vector(7 downto 0);
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        en              : in     vl_logic;
        up              : in     vl_logic
    );
end Counter_10927143;
