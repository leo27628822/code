library verilog;
use verilog.vl_types.all;
entity TM_AddSub4 is
end TM_AddSub4;
