library verilog;
use verilog.vl_types.all;
entity tb_Pipelined is
end tb_Pipelined;
