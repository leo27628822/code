library verilog;
use verilog.vl_types.all;
entity TM_RCA4 is
end TM_RCA4;
