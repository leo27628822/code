library verilog;
use verilog.vl_types.all;
entity stimulus is
end stimulus;
