library verilog;
use verilog.vl_types.all;
entity Simulate is
end Simulate;
