library verilog;
use verilog.vl_types.all;
entity simulate is
end simulate;
