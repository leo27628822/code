library verilog;
use verilog.vl_types.all;
entity Stimulate is
end Stimulate;
